module included();
endmodule
