module included();
endmodule
module include();
endmodule
