`include "./included.v"

module include();
endmodule
